`timescale 1ns/1ps
module xor1(a,b,c);
input a,b;
output c;
assign c = (a^b);
endmodule